
--******************************************************--
--        PONTIFICIA UNIVERSIDAD JAVERIANA              --
--                Disegno Digital                       --
--          Seccion de Tecnicas Digitales               --
-- 													              --
-- Titulo :                                             --
-- Fecha  :  	D:XX M:XX Y:20XX                         --
--******************************************************--

LIBRARY IEEE;
USE IEEE.std_logic_1164.all;
LIBRARY ALTERA;
USE ALTERA.altera_primitives_components.all;

--******************************************************--
-- Comentarios:
-- 
-- 
--******************************************************--

ENTITY StateTransform IS
	
	PORT	 (
				Qs    : IN  STD_LOGIC_VECTOR(85 DOWNTO 0);
				State : OUT STD_LOGIC_VECTOR( 6 DOWNTO 0)
			 );
	
END ENTITY StateTransform;

ARCHITECTURE StateTransformArch OF StateTransform IS

BEGIN

--******************************************************--
-- 
-- 
-- 
--******************************************************--

WITH Qs SELECT
State <= "0000000" WHEN "00000000000000000000000000000000000000000000000000000000000000000000000000000000000001",
         "0000001" WHEN "00000000000000000000000000000000000000000000000000000000000000000000000000000000000010",
			"0000010" WHEN "00000000000000000000000000000000000000000000000000000000000000000000000000000000000100",
			"0000011" WHEN "00000000000000000000000000000000000000000000000000000000000000000000000000000000001000",
			"0000100" WHEN "00000000000000000000000000000000000000000000000000000000000000000000000000000000010000",
			"0000101" WHEN "00000000000000000000000000000000000000000000000000000000000000000000000000000000100000",
			"0000110" WHEN "00000000000000000000000000000000000000000000000000000000000000000000000000000001000000",
			"0000111" WHEN "00000000000000000000000000000000000000000000000000000000000000000000000000000010000000",
			"0001000" WHEN "00000000000000000000000000000000000000000000000000000000000000000000000000000100000000",
			"0001001" WHEN "00000000000000000000000000000000000000000000000000000000000000000000000000001000000000",
			"0001010" WHEN "00000000000000000000000000000000000000000000000000000000000000000000000000010000000000",
			"0001011" WHEN "00000000000000000000000000000000000000000000000000000000000000000000000000100000000000",
			"0001100" WHEN "00000000000000000000000000000000000000000000000000000000000000000000000001000000000000",
			"0001101" WHEN "00000000000000000000000000000000000000000000000000000000000000000000000010000000000000",
			"0001110" WHEN "00000000000000000000000000000000000000000000000000000000000000000000000100000000000000",
			"0001111" WHEN "00000000000000000000000000000000000000000000000000000000000000000000001000000000000000",
			"0010000" WHEN "00000000000000000000000000000000000000000000000000000000000000000000010000000000000000",
			"0010001" WHEN "00000000000000000000000000000000000000000000000000000000000000000000100000000000000000",
			"0010010" WHEN "00000000000000000000000000000000000000000000000000000000000000000001000000000000000000",
			"0010011" WHEN "00000000000000000000000000000000000000000000000000000000000000000010000000000000000000",
			"0010100" WHEN "00000000000000000000000000000000000000000000000000000000000000000100000000000000000000",
			"0010101" WHEN "00000000000000000000000000000000000000000000000000000000000000001000000000000000000000",
			"0010110" WHEN "00000000000000000000000000000000000000000000000000000000000000010000000000000000000000",
			"0010111" WHEN "00000000000000000000000000000000000000000000000000000000000000100000000000000000000000",
			"0011000" WHEN "00000000000000000000000000000000000000000000000000000000000001000000000000000000000000",
			"0011001" WHEN "00000000000000000000000000000000000000000000000000000000000010000000000000000000000000",
			"0011010" WHEN "00000000000000000000000000000000000000000000000000000000000100000000000000000000000000",
			"0011011" WHEN "00000000000000000000000000000000000000000000000000000000001000000000000000000000000000",
			"0011100" WHEN "00000000000000000000000000000000000000000000000000000000010000000000000000000000000000",
			"0011101" WHEN "00000000000000000000000000000000000000000000000000000000100000000000000000000000000000",
			"0011110" WHEN "00000000000000000000000000000000000000000000000000000001000000000000000000000000000000",
			"0011111" WHEN "00000000000000000000000000000000000000000000000000000010000000000000000000000000000000",
			"0100000" WHEN "00000000000000000000000000000000000000000000000000000100000000000000000000000000000000",
			"0100001" WHEN "00000000000000000000000000000000000000000000000000001000000000000000000000000000000000",
			"0100010" WHEN "00000000000000000000000000000000000000000000000000010000000000000000000000000000000000",
			"0100011" WHEN "00000000000000000000000000000000000000000000000000100000000000000000000000000000000000",
			"0100100" WHEN "00000000000000000000000000000000000000000000000001000000000000000000000000000000000000",
			"0100101" WHEN "00000000000000000000000000000000000000000000000010000000000000000000000000000000000000",
			"0100110" WHEN "00000000000000000000000000000000000000000000000100000000000000000000000000000000000000",
			"0100111" WHEN "00000000000000000000000000000000000000000000001000000000000000000000000000000000000000",
			"0101000" WHEN "00000000000000000000000000000000000000000000010000000000000000000000000000000000000000",
			"0101001" WHEN "00000000000000000000000000000000000000000000100000000000000000000000000000000000000000",
			"0101010" WHEN "00000000000000000000000000000000000000000001000000000000000000000000000000000000000000",
			"0101011" WHEN "00000000000000000000000000000000000000000010000000000000000000000000000000000000000000",
			"0101100" WHEN "00000000000000000000000000000000000000000100000000000000000000000000000000000000000000",
			"0101101" WHEN "00000000000000000000000000000000000000001000000000000000000000000000000000000000000000",
			"0101110" WHEN "00000000000000000000000000000000000000010000000000000000000000000000000000000000000000",
			"0101111" WHEN "00000000000000000000000000000000000000100000000000000000000000000000000000000000000000",
			"0110000" WHEN "00000000000000000000000000000000000001000000000000000000000000000000000000000000000000",
			"0110001" WHEN "00000000000000000000000000000000000010000000000000000000000000000000000000000000000000",
			"0110010" WHEN "00000000000000000000000000000000000100000000000000000000000000000000000000000000000000",
			"0110011" WHEN "00000000000000000000000000000000001000000000000000000000000000000000000000000000000000",
			"0110100" WHEN "00000000000000000000000000000000010000000000000000000000000000000000000000000000000000",
			"0110101" WHEN "00000000000000000000000000000000100000000000000000000000000000000000000000000000000000",
			"0110110" WHEN "00000000000000000000000000000001000000000000000000000000000000000000000000000000000000",
			"0110111" WHEN "00000000000000000000000000000010000000000000000000000000000000000000000000000000000000",
			"0111000" WHEN "00000000000000000000000000000100000000000000000000000000000000000000000000000000000000",
			"0111001" WHEN "00000000000000000000000000001000000000000000000000000000000000000000000000000000000000",
			"0111010" WHEN "00000000000000000000000000010000000000000000000000000000000000000000000000000000000000",
			"0111011" WHEN "00000000000000000000000000100000000000000000000000000000000000000000000000000000000000",
			"0111100" WHEN "00000000000000000000000001000000000000000000000000000000000000000000000000000000000000",
			"0111101" WHEN "00000000000000000000000010000000000000000000000000000000000000000000000000000000000000",
			"0111110" WHEN "00000000000000000000000100000000000000000000000000000000000000000000000000000000000000",
			"0111111" WHEN "00000000000000000000001000000000000000000000000000000000000000000000000000000000000000",
			"1000001" WHEN "00000000000000000000010000000000000000000000000000000000000000000000000000000000000000",
			"1000010" WHEN "00000000000000000000100000000000000000000000000000000000000000000000000000000000000000",
			"1000011" WHEN "00000000000000000001000000000000000000000000000000000000000000000000000000000000000000",
			"1000100" WHEN "00000000000000000010000000000000000000000000000000000000000000000000000000000000000000",
			"1000101" WHEN "00000000000000000100000000000000000000000000000000000000000000000000000000000000000000",
			"1000110" WHEN "00000000000000001000000000000000000000000000000000000000000000000000000000000000000000",
			"1000111" WHEN "00000000000000010000000000000000000000000000000000000000000000000000000000000000000000",
			"1001000" WHEN "00000000000000100000000000000000000000000000000000000000000000000000000000000000000000",
			"1001001" WHEN "00000000000001000000000000000000000000000000000000000000000000000000000000000000000000",
			"1001010" WHEN "00000000000010000000000000000000000000000000000000000000000000000000000000000000000000",
			"1001011" WHEN "00000000000100000000000000000000000000000000000000000000000000000000000000000000000000",
			"1001100" WHEN "00000000001000000000000000000000000000000000000000000000000000000000000000000000000000",
			"1001101" WHEN "00000000010000000000000000000000000000000000000000000000000000000000000000000000000000",
			"1001110" WHEN "00000000100000000000000000000000000000000000000000000000000000000000000000000000000000",
			"1001111" WHEN "00000001000000000000000000000000000000000000000000000000000000000000000000000000000000",
			"1010000" WHEN "00000010000000000000000000000000000000000000000000000000000000000000000000000000000000",
			"1010001" WHEN "00000100000000000000000000000000000000000000000000000000000000000000000000000000000000",
			"1010010" WHEN "00001000000000000000000000000000000000000000000000000000000000000000000000000000000000",
			"1010011" WHEN "00010000000000000000000000000000000000000000000000000000000000000000000000000000000000",
			"1010100" WHEN "00100000000000000000000000000000000000000000000000000000000000000000000000000000000000",
			"1010101" WHEN "01000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
			"1010110" WHEN "10000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
			"1111110" WHEN "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
			"1111111" WHEN OTHERS;

--******************************************************--
-- 
-- Summon This Block:
-- 
--******************************************************--
--BlockN: ENTITY WORK.StateTransform 
--PORT MAP	  (Qs    => SLV,
--				State => SLV
--			  );
--******************************************************--

END StateTransformArch;